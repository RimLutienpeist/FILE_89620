`timescale 1ns / 1ps

module Mux4to1b4_tb;


  reg  [1:0] S;
  reg  [3:0] D0, D1, D2, D3;

  wire [3:0] Y;

  Mux4to1b4 uut (
    .S(S),
    .D0(D0),
    .D1(D1),
    .D2(D2),
    .D3(D3),
    .Y(Y)
  );

  initial begin
  for (S = 0; ; S = S + 1) begin
    case(S)
      2'b00: begin
        D0 = 4'b1111;
        D1 = 4'b0000;
        D2 = 4'b0000;
        D3 = 4'b0000;
        #5;  
        D0 = 4'b1010;
        D1 = 4'b0101;
        D2 = 4'b1100;
        D3 = 4'b0011;
        #5;  
        D0 = 4'b1111;
        D1 = 4'b1111;
        D2 = 4'b0000;
        D3 = 4'b0000;
        #5;
        D0 = 4'b1100;
        D1 = 4'b0110;
        D2 = 4'b0011;
        D3 = 4'b1001;
      end
      2'b01: begin
        D0 = 4'b1111;
        D1 = 4'b0000;
        D2 = 4'b0000;
        D3 = 4'b0000;
        #5;  
        D0 = 4'b1010;
        D1 = 4'b0101;
        D2 = 4'b1100;
        D3 = 4'b0011;
        #5;  
        D0 = 4'b1111;
        D1 = 4'b1111;
        D2 = 4'b0000;
        D3 = 4'b0000;
        #5;
        D0 = 4'b1100;
        D1 = 4'b0110;
        D2 = 4'b0011;
        D3 = 4'b1001;
      end
      2'b10: begin
        D0 = 4'b1111;
        D1 = 4'b0000;
        D2 = 4'b0000;
        D3 = 4'b0000;
        #5;  
        D0 = 4'b1010;
        D1 = 4'b0101;
        D2 = 4'b1100;
        D3 = 4'b0011;
        #5;  
        D0 = 4'b1111;
        D1 = 4'b1111;
        D2 = 4'b0000;
        D3 = 4'b0000;
        #5;
        D0 = 4'b1100;
        D1 = 4'b0110;
        D2 = 4'b0011;
        D3 = 4'b1001;
      end
      2'b11: begin
        D0 = 4'b1111;
        D1 = 4'b0000;
        D2 = 4'b0000;
        D3 = 4'b0000;
        #5;  
        D0 = 4'b1010;
        D1 = 4'b0101;
        D2 = 4'b1100;
        D3 = 4'b0011;
        #5;  
        D0 = 4'b1111;
        D1 = 4'b1111;
        D2 = 4'b0000;
        D3 = 4'b0000;
        #5;
        D0 = 4'b1100;
        D1 = 4'b0110;
        D2 = 4'b0011;
        D3 = 4'b1001;
        #10
        $finish;
      end
    endcase
    #10;  
    end
  end

endmodule